----------------------------------------------------------------------------------
-- Compa��a:            Estado Finito
-- Ingeniero:           Carlos Ramos
-- 
-- Fecha de creaci�n:   2013/06/01 19:23:01
-- Nombre del m�dulo:   contador_servo_pwm - Behavioral
-- Descripci�n: 
--   Contador de 0 a 127, cuyo valor incrementa o decrementa gracias a un bot�n
--   para cada funci�n (un bot�n incrementa, un bot�n decrementa).
--
-- Comentarios adicionales:
--   Se puede encontrar m�s informaci�n en la siguiente direcci�n:
--   http://www.estadofinito.com/control-servomotor-dos-botones/
--
-- Revisi�n:
--   Revisi�n 0.01 - Archivo creado.
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity contador_servo_pwm is
    PORT (
        clk   : IN  STD_LOGIC; -- Reloj de 64kHz.
        reset : IN  STD_LOGIC; -- Bot�n de reset.
		cnt_up: IN  STD_LOGIC; -- Bot�n de incremento.
		cnt_dn: IN  STD_LOGIC; -- Bot�n de decremento.
        pos   : OUT STD_LOGIC_VECTOR(6 downto 0) -- Salida a servomotor.
    );
end contador_servo_pwm;

architecture Behavioral of contador_servo_pwm is
	-- Se�al utilizada para modificar la salida "pos".
	signal contador: UNSIGNED(6 downto 0) := (OTHERS => '0');
begin
	proceso_contador: process (clk, reset, cnt_up, cnt_dn) begin
		if (reset = '1') then
			contador <= (others => '0');
		elsif rising_edge(clk) then
			if (cnt_up = '1' AND contador < 127) then
				contador <= contador + 1;
			elsif (cnt_dn = '1' AND contador > 0) then
				contador <= contador - 1;
			end if;
		end if;
	end process;
	
	-- Asignaci�n del valor del contador a la salida del m�dulo.
	pos <= STD_LOGIC_VECTOR(contador);
end Behavioral;